module cond_unit ()


endmodule